module ysyx_23060240_SRAM_LSU(
    input clk,

)
endmodule